// Tutorial 5 Parte 2 - Register bank
//
module register_bank #(
   parameter WIDTH = 8 )
 (
   input                   clk,
   input                   rst,
   input                   wr_en,
   input       [WIDTH-1:0] in,
   output      [WIDTH-1:0] out
);
   

endmodule
