// Tutorial 1 - 1 bit full adder
//
module onebitadder (
  input a, b, cin,
  output sum, cout
);

endmodule
