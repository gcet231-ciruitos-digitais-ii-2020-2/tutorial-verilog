// Tutorial 6 - Datapath completo.

module top #(
   parameter WIDTH = 8
   )(
   input clk,
   input rst,
   input [5:0] cmdin,
   input [WIDTH-1:0] din_1,
   input [WIDTH-1:0] din_2,
   input [WIDTH-1:0] din_3,
   output [WIDTH-1:0] dout_low,
   output [WIDTH-1:0] dout_high,
   output zero,
   output error
);


endmodule
