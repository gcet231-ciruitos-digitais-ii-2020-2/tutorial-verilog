// Tutorial 5 Parte 1 - Parameterized 4-input MUX
//
module mux4 #( 
  parameter WIDTH = 8
  )(
  input      [WIDTH-1:0] din1, din2, din3, din4,
  input      [1:0]       select,     
  output     [WIDTH-1:0] dout 
);


endmodule
