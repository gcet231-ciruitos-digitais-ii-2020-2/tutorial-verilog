// Tutorial 5 Parte 3 - Basic ALU

module alu #(
   parameter WIDTH = 8
   )(
   input [WIDTH-1:0]    in1, in2,
   input [3:0]          op,
   input nvalid_data,
   output [2*WIDTH-1:0]  out,
   output  zero, 
   output error
);


endmodule
